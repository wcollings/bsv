aaaa,b,c,d1.000000e+00�2.000000e+00�3.000000e+00�4.000000e+00�5.000000e+00�6.000000e+00�7.000000e+00�8.000000e+00�8.000000e+00�